/* Unidade multiplicadora (MUU - MUltiplication Unit):
 *	Realiza operacoes relacionadas a multiplicacao e divisao. Guarda os
 * resultados nos registradores 'hi' e 'lo', que devem ser resgatados posterior-
 * mente, dependendo da operacao.
 */
/*----------------------------------------------------------------------------*/
module multiplilcation_unit (
	input [31:0] rs, rt,		// Operandos
	input [3:0] operation,	// Operacao - pode ser reduzido p/ 3 bits,
									// deixando 4 para eventual expansao
	output div_zero,			// Indica divisao por zero
	output reg [31:0] out,	// Saida para os 32 bits SUPERIORES [63:32]
	);
	
	reg [63:0] result;
	reg [31:0] hi, lo;
	
	always @(*) begin
		div_zero <= 0;
		
		case(operation)
			4'b0000: begin	// MUL
				result <= $signed(rs) * $signed(rt);
				out <= result[31:0];
			end
			
			4'b0001: begin	// MULT
				result <= $signed(rs) * $signed(rt);
				hi <= result[64:32];
				lo <= result[31:0];
			end
			
			4'b0010: begin	// MADD
				result <= $signed(rs) * $signed(rt);
				hi <= hi + result[64:32];
				lo <= lo + result[31:0];
			end
			
			4'b0011: begin	// MSUBU: multip., neste caso, desconsidera sinal
				result <= rs * rt;
				hi <= hi - result[64:32];
				lo <= lo - result[31:0];
			end
			
			4'b0100: begin // DIV
				if (B != 0) begin
					lo <= $signed(A) / $signed(B);
					hi <= $signed(A) % $signed(B);
				end
				
				else begin
					div_zero = 1'b1;
				end
				
			4'b0101:	// MFHI
				out <= hi;
			end
			
			4'b0110:	// MFLO
				out <= lo;
			end
			
		endcase
	end
	
endmodule